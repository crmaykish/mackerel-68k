module system_controller(
	input RST_n,
	input CLK_n
);



endmodule
